// Here, and_gate is user defined module name
// "a", "b", "out" are userdefined pandt names
module and_gate (a, b, out);
input a, b;
output out;
// "and" is a data type for creating data type
and and1(out, a, b);
endmodule